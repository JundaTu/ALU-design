library ieee;
library work;
use ieee.std_logic_1164.all;
use work.add_sub_32;

entity add_sub_32_test is
  
end add_sub_32_test;

architecture behavior of add_sub_32_test is
signal a,b,sum : std_logic_vector(31 downto 0);
signal cout,invert: std_logic;

component add_sub_32 is
  port(
    a : in std_logic_vector(31 downto 0);
    b : in std_logic_vector(31 downto 0);
    invert : in std_logic;
    cout : out std_logic;
    sum : out std_logic_vector(31 downto 0)
  );
end component add_sub_32;

begin
  test_comp : add_sub_32
  port map(
  a=>a,
  b=>b,
  invert=>invert,
  cout=>cout,
  sum=>sum
  );
  testbench : process
  begin
    invert<='0';
    a<="00000000000000000000000000000000";
    b<="00000000000000000000000000000000";
    
    wait for 50 ns;
    a<="00000000000000000000000000000001";
    b<="00000000000000000000000000000000";
    wait for 50ns;
    wait for 50 ns;
    a<="00000000000000000000000000000001";
    b<="00000000000000000000000000000001";
    wait for 50 ns;
    a<="00000000000000000000000000000001";
    b<="00000000000000000000000000000010";
    wait for 50 ns;
    a<="00000000000000000000000000000001";
    b<="01111111111111111111111111111111";
    wait for 50 ns;
    a<="00000000000000000000000000000001";
    b<="11111111111111111111111111111111";
    wait for 50 ns;
    a<="11111111111111111111111111111111";
    b<="00000000000000000000000000000111";
    invert<='1';
    wait;
    
  end process;
end architecture behavior;








